import Vector::*;

typedef 80 InstSz;
typedef Bit#(InstSz) Inst; 

typedef 64 AddrSz;
typedef Bit#(AddrSz) Addr;

typedef 64 DataSz;
typedef Bit#(DataSz) Data;

typedef Bit#(8) Byte;



